module hello();
  
	initial begin //usa quando está descrevendo o testebanch
		$display("*** Hello World ***"); //imprime string na tela
      
    $finish(); //para a simulação
      
	end
  
endmodule: hello;
